[aimspice]
[description]
475
TG Switch

.include gpdk90nm_tt.cir

.param lp = 1U
.param wp = 1U
.param ln = 1U
.param wn = 1U


Vdd1 1 0 dc 0
Vdd2 4 0 dc 1
VPULSE1 2 0 PULSE(0 1 0 1ns 1ns 50ns 200ns)
*VPULSE2 1 0 PULSE(0 1 0 1ns 1ns 50ns 100ns)
*VPULSE3 4 0 PULSE(1 0 0 1ns 1ns 50ns 100ns)
	
*XMN1 6 5 0 0 nmos1v L=ln W=wn
*XMP1 6 5 1 1 pmos1v L=lp W=wp
*d g s b
XMP2 2 1 3 3 pmos1v L=lp W=wp
XMN2 2 4 3 3 nmos1v L=lp W=wn
C1 3 0 100fF

.plot tran V(2) V(3)
.plot tran V(1) V(4)

[tran]
1ns
500ns
X
X
0
[ana]
4 0
[end]
