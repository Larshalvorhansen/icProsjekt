[aimspice]
[description]
453
NOR GATE

.include gpdk90nm_tt.cir

.param LP = 0.1U
.param WP = 1U
.param LN = 0.1U
.param WN = 1U

.subckt NOR in1 in2 out vdd GND
XMP1 2 in1 vdd vdd PMOS1V L=LP W=WP
XMP2 out in2 2 vdd PMOS1V L=LP W=WP
XMN1 out in1 GND GND NMOS1V L=LN W=WN
XMN2 out in2 GND GND NMOS1V L=LN W=WN
.ends

vdd1 1 0 dc 1
VPULSE 2 0 PULSE(0 1 0 40ns 1ns 1ns 100ns)
vin2 3 0 PULSE(0 1 0 40ns 1ns 1ns 150ns)

XNOR1 2 3 4 1 0 NOR
.plot tran V(2) V(3) V(4)
[tran]
1ns
500ns
X
X
0
[ana]
4 0
[end]
