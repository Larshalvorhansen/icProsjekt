[aimspice]
[description]
555
AND GATE2

.include gpdk90nm_tt.cir

.param LP = 0.1U
.param WP = 1U
.param LN = 0.1U
.param WN = 1U
*d g s b
.subckt AND in1 in2 out VDD GND
XMN1 out in1 GND GND nmos1V L=LN W=WN
XMN2 out in2 GND GND nmos1V L=LN W=WN
XMP1 1 in1 VDD VDD nmos1V L=LP W=WP
XMP2 out in2 1 1 nmos1V L=LP W=WP
.ends

*PULSE Initial value Pulsed value Delay time Rise time Fall time Pulse width Period
vdd1 1 0 dc 1
VPULSE 2 0 PULSE(0 1 0 1ns 1ns 50ns 100ns)
vin2 3 0 PULSE(0 1 0 1ns 1ns 75ns 150ns)

XAND1 2 3 4 1 0 AND
.plot tran V(2) V(3) V(4)





[tran]
1ns
500ns
X
X
0
[ana]
4 0
[end]
