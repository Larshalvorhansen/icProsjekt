[aimspice]
[description]
300
NOR GATE

.include gpdk90nm_tt.cir

.param lp = 0.1U
.param wp = 1U
.param ln = 0.1U
.param wn = 1U

.subckt NOR vdd GND in1 in2 out:
XMP1 2 in1 vdd vdd PMOS1V L=LP W=WP
XMP2 out in2 2 vdd PMOS1V L=LP W=WP
XMN1 out in1 GND GND NMOS1V L=LN W=WN
XMN2 out in2 GND GND NMOS1V L=LN W=WN



[end]
