[aimspice]
[description]
470
AND GATE2

.include gpdk90nm_tt.cir

.param LP = 0.1U
.param WP = 1U
.param LN = 0.1U
.param WN = 1U
*d g s b

XMN1 2 3 1 1 nmos1V L=LN W=WN
XMN2 5 4 2 2 nmos1V L=LN W=WN
XMP1 5 3 0 0 nmos1V L=LP W=WP
XMP2 5 4 0 0 nmos1V L=LP W=WP


*PULSE Initial value Pulsed value Delay time Rise time Fall time Pulse width Period
vdd1 1 0 dc 1
vin1 3 0 PULSE(0 1 0 1ns 1ns 50ns 100ns)
vin2 4 0 PULSE(0 1 0 1ns 1ns 50ns 200ns)

.plot tran V(5) V(3) V(4)





[tran]
1ns
500ns
X
X
0
[ana]
4 0
[end]
