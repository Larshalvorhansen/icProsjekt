[aimspice]
[description]
305
TG Switch
Vdd1 1 0 dc 0 
Vdd2 4 0 dc 5

.include gpdk90nm_tt.cir

.param LP = 1U
.param WP = 1U
.param LN = 1U
.param WN = 1U

VPULSE 2 0 PULSE 0 1 0S 0US 50US 100US

XMP1 2 1 3 3 PMOS1V L=LP W=WP
XMN1 2 4 3 3 NMOS1V L=LN W=WN 
C1 3 0 100fF

.plot tran V(2) !5.2
.plot tran V(3) !5.2


[dc]
1
vin
0
1
0.01
[tran]
1ns
100ns
X
X
0
[ana]
4 0
[end]
