[aimspice]
[description]
294
AND GATE

.include gpdk90nm_tt.cir

.param lp = 0.1U
.param wp = 1U
.param ln = 0.1U
.param wn = 1U

.subckt AND vdd GND in1 in2 out:
XMP1 GND in1 out vdd PMOS1V L=LP W=WP
XMP2 GND in2 out vdd PMOS1V L=LP W=WP
XMN1 vdd in1 3 GND NMOS1V L=LN W=WN
XMN2 3 in2 out GND NMOS1V L=LN W=WN
[end]
