[aimspice]
[description]
305
TG Switch
Vdd1 1 0 dc 0


.include gpdk90nm_tt.cir
.include Inverter.cir

.param LP = 1U
.param WP = 1U
.param LN = 1U
.param WN = 1U

VPULSE 2 0 PULSE 0 1 0S 0US 50US 100US

*d g s b
XMP1 1 5 2 1 PMOS1V L=LP W=WP
XMN1 2 6 1 0 NMOS1V L=LN W=WN
Xinv 1 0 5 6 invert
*vdd vss in out

.plot tran V(2) 
.plot tran V(3)