[aimspice]
[description]
242
Inverter Subcircuit

.include gpdk90nm_tt.cir
.param lp = 0.1U
.param wp = 1U
.param ln = 0.1U
.param wn = 1U



.subckt invert in out vdd vss 
XMN1 out in vss vss nmos1v L=ln W=wn
XMP1 out in vdd vdd pmos1v L=lp W=wp
.ends



[dc]
1
vin
0
1
0.01
[ana]
1 0
[end]
